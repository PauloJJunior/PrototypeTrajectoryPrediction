{"lastScore":0,"coins":0,"currentLevel":1,"rounds":0,"currentCharacter":0,"maxLevel":4}