{"coins":7,"currentLevel":3,"playerMaxLevel":1,"maxLevel":1}