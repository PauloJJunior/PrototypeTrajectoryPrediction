{"coins":4,"currentLevel":3,"playerMaxLevel":1,"maxLevel":1}